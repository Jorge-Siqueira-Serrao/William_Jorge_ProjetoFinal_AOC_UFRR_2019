LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY memoria_ram IS
    PORT (
        clock : IN std_logic;
        mem_write : IN std_logic;
        mem_read : IN std_logic;
        endereco : IN std_logic_vector(7 DOWNTO 0);
        in_port : IN std_logic_vector(7 DOWNTO 0);
        out_port : OUT std_logic_vector(7 DOWNTO 0)
    );
END memoria_ram;

ARCHITECTURE behavior OF memoria_ram IS
    TYPE memoriaRam IS ARRAY (0 TO 7) OF std_logic_vector(7 DOWNTO 0);
    SIGNAL ram : memoriaRam := (OTHERS => "00000000");
BEGIN
    PROCESS (clock)
    BEGIN
        IF rising_edge(clock) THEN
            IF (mem_write = '1') THEN
                ram(to_integer(unsigned(endereco))) <= in_port;
            END IF;
            IF (mem_read = '1') THEN
                out_port <= ram(to_integer(unsigned(endereco)));
            END IF;
        END IF;
    END PROCESS;
END behavior;